library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity vc707_prom_flasher is
--  Port ( );
end vc707_prom_flasher;

architecture Behavioral of vc707_prom_flasher is

begin


end Behavioral;
