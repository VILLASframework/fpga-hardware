`timescale 1ns / 1ps

/* Macro definitions.
 *
 * @author Hatim Kanchwala <hatim@hatimak.me>
 * @copyright 2019 Hatim Kanchwala
 */

`ifndef DEFINES_VH
 `define DEFINES_VH

`endif
