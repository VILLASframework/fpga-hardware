`timescale 1ns / 1ps

/* Macro definitions.
 *
 * @author Hatim Kanchwala <hatim@hatimak.me>
 * @copyright 2019 Hatim Kanchwala
 */

// `define INCLUDE_ILA_AURORA_PRE
`define INCLUDE_ILA_AURORA
// `define INCLUDE_ILA_AURORA_POST
